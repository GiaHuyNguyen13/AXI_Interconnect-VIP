module tb;
  reg clk;
  
  always #10 clk =~ clk;
  interface _if (clk);

  
  initial begin
    clk <= 0;
    uvm_config_db#(virtual interface)::set(null, "uvm_test_top", "interface", _if);
    run_test("");
  end

  initial begin
    $vcdplusfile("wave_wave.vpd");
    $vcdpluson();
  end

  // Instantiate DUT
  axi_interconnect_wrap_2x2 dut(
    .clk (clk),
    .rst (rst),

    /*
     * AXI slave interface
     */
    .s00_axi_awid (_if.s00_axi_awid),
    .s00_axi_awaddr (_if.s00_axi_awaddr),
    .s00_axi_awlen (_if.s00_axi_awlen),
    .s00_axi_awsize (_if.s00_axi_awsize),
    .s00_axi_awburst (_if.s00_axi_awburst),
    .s00_axi_awlock (_if.s00_axi_awlock),
    .s00_axi_awcache (_if.s00_axi_awcache),
    .s00_axi_awprot (_if.s00_axi_awprot),
    .s00_axi_awqos (_if.s00_axi_awqos),
    .s00_axi_awuser (_if.s00_axi_awuser),
    .s00_axi_awvalid (_if.s00_axi_awvalid),
    .s00_axi_awready (_if.s00_axi_awready),
    .s00_axi_wdata (_if.s00_axi_wdata),
    .s00_axi_wstrb (_if.s00_axi_wstrb),
    .s00_axi_wlast (_if.s00_axi_wlast),
    .s00_axi_wuser (_if.s00_axi_wuser),
    .s00_axi_wvalid (_if.s00_axi_wvalid),
    .s00_axi_wready (_if.s00_axi_wready),
    .s00_axi_bid (_if.s00_axi_bid),
    .s00_axi_bresp (_if.s00_axi_bresp),
    .s00_axi_buser (_if.s00_axi_buser),
    .s00_axi_bvalid (_if.s00_axi_bvalid),
    .s00_axi_bready (_if.s00_axi_bready),
    .s00_axi_arid (_if.s00_axi_arid),
    .s00_axi_araddr (_if.s00_axi_araddr),
    .s00_axi_arlen (_if.s00_axi_arlen),
    .s00_axi_arsize (_if.s00_axi_arsize),
    .s00_axi_arburst (_if.s00_axi_arburst),
    .s00_axi_arlock (_if.s00_axi_arlock),
    .s00_axi_arcache (_if.s00_axi_arcache),
    .s00_axi_arprot (_if.s00_axi_arprot),
    .s00_axi_arqos (_if.s00_axi_arqos),
    .s00_axi_aruser (_if.s00_axi_aruser),
    .s00_axi_arvalid (_if.s00_axi_arvalid),
    .s00_axi_arready (_if.s00_axi_arready),
    .s00_axi_rid (_if.s00_axi_rid),
    .s00_axi_rdata (_if.s00_axi_rdata),
    .s00_axi_rresp (_if.s00_axi_rresp),
    .s00_axi_rlast (_if.s00_axi_rlast),
    .s00_axi_ruser (_if.s00_axi_ruser),
    .s00_axi_rvalid (_if.s00_axi_rvalid),
    .s00_axi_rready (_if.s00_axi_rready),

    .s01_axi_awid (_if.s01_axi_awid),
    .s01_axi_awaddr (_if.s01_axi_awaddr),
    .s01_axi_awlen (_if.s01_axi_awlen),
    .s01_axi_awsize (_if.s01_axi_awsize),
    .s01_axi_awburst (_if.s01_axi_awburst),
    .s01_axi_awlock (_if.s01_axi_awlock),
    .s01_axi_awcache (_if.s01_axi_awcache),
    .s01_axi_awprot (_if.s01_axi_awprot),
    .s01_axi_awqos (_if.s01_axi_awqos),
    .s01_axi_awuser (_if.s01_axi_awuser),
    .s01_axi_awvalid (_if.s01_axi_awvalid),
    .s01_axi_awready (_if.s01_axi_awready),
    .s01_axi_wdata (_if.s01_axi_wdata),
    .s01_axi_wstrb (_if.s01_axi_wstrb),
    .s01_axi_wlast (_if.s01_axi_wlast),
    .s01_axi_wuser (_if.s01_axi_wuser),
    .s01_axi_wvalid (_if.s01_axi_wvalid),
    .s01_axi_wready (_if.s01_axi_wready),
    .s01_axi_bid (_if.s01_axi_bid),
    .s01_axi_bresp (_if.s01_axi_bresp),
    .s01_axi_buser (_if.s01_axi_buser),
    .s01_axi_bvalid (_if.s01_axi_bvalid),
    .s01_axi_bready (_if.s01_axi_bready),
    .s01_axi_arid (_if.s01_axi_arid),
    .s01_axi_araddr (_if.s01_axi_araddr),
    .s01_axi_arlen (_if.s01_axi_arlen),
    .s01_axi_arsize (_if.s01_axi_arsize),
    .s01_axi_arburst (_if.s01_axi_arburst),
    .s01_axi_arlock (_if.s01_axi_arlock),
    .s01_axi_arcache (_if.s01_axi_arcache),
    .s01_axi_arprot (_if.s01_axi_arprot),
    .s01_axi_arqos (_if.s01_axi_arqos),
    .s01_axi_aruser (_if.s01_axi_aruser),
    .s01_axi_arvalid (_if.s01_axi_arvalid),
    .s01_axi_arready (_if.s01_axi_arready),
    .s01_axi_rid (_if.s01_axi_rid),
    .s01_axi_rdata (_if.s01_axi_rdata),
    .s01_axi_rresp (_if.s01_axi_rresp),
    .s01_axi_rlast (_if.s01_axi_rlast),
    .s01_axi_ruser (_if.s01_axi_ruser),
    .s01_axi_rvalid (_if.s01_axi_rvalid),
    .s01_axi_rready (_if.s01_axi_rready),

    /*
     * AXI master interface
     */
    .m00_axi_awid (_if.m00_axi_awid),
    .m00_axi_awaddr (_if.m00_axi_awaddr),
    .m00_axi_awlen (_if.m00_axi_awlen),
    .m00_axi_awsize (_if.m00_axi_awsize),
    .m00_axi_awburst (_if.m00_axi_awburst),
    .m00_axi_awlock (_if.m00_axi_awlock),
    .m00_axi_awcache (_if.m00_axi_awcache),
    .m00_axi_awprot (_if.m00_axi_awprot),
    .m00_axi_awqos (_if.m00_axi_awqos),
    .m00_axi_awregion (_if.m00_axi_awregion),
    .m00_axi_awuser (_if.m00_axi_awuser),
    .m00_axi_awvalid (_if.m00_axi_awvalid),
    .m00_axi_awready (_if.m00_axi_awready),
    .m00_axi_wdata (_if.m00_axi_wdata),
    .m00_axi_wstrb (_if.m00_axi_wstrb),
    .m00_axi_wlast (_if.m00_axi_wlast),
    .m00_axi_wuser (_if.m00_axi_wuser),
    .m00_axi_wvalid (_if.m00_axi_wvalid),
    .m00_axi_wready (_if.m00_axi_wready),
    .m00_axi_bid (_if.m00_axi_bid),
    .m00_axi_bresp (_if.m00_axi_bresp),
    .m00_axi_buser (_if.m00_axi_buser),
    .m00_axi_bvalid (_if.m00_axi_bvalid),
    .m00_axi_bready (_if.m00_axi_bready),
    .m00_axi_arid (_if.m00_axi_arid),
    .m00_axi_araddr (_if.m00_axi_araddr),
    .m00_axi_arlen (_if.m00_axi_arlen),
    .m00_axi_arsize (_if.m00_axi_arsize),
    .m00_axi_arburst (_if.m00_axi_arburst),
    .m00_axi_arlock (_if.m00_axi_arlock),
    .m00_axi_arcache (_if.m00_axi_arcache),
    .m00_axi_arprot (_if.m00_axi_arprot),
    .m00_axi_arqos (_if.m00_axi_arqos),
    .m00_axi_arregion (_if.m00_axi_arregion),
    .m00_axi_aruser (_if.m00_axi_aruser),
    .m00_axi_arvalid (_if.m00_axi_arvalid),
    .m00_axi_arready (_if.m00_axi_arready),
    .m00_axi_rid (_if.m00_axi_rid),
    .m00_axi_rdata (_if.m00_axi_rdata),
    .m00_axi_rresp (_if.m00_axi_rresp),
    .m00_axi_rlast (_if.m00_axi_rlast),
    .m00_axi_ruser (_if.m00_axi_ruser),
    .m00_axi_rvalid (_if.m00_axi_rvalid),
    .m00_axi_rready (_if.m00_axi_rready),

    .m01_axi_awid (_if.m01_axi_awid),
    .m01_axi_awaddr (_if.m01_axi_awaddr),
    .m01_axi_awlen (_if.m01_axi_awlen),
    .m01_axi_awsize (_if.m01_axi_awsize),
    .m01_axi_awburst (_if.m01_axi_awburst),
    .m01_axi_awlock (_if.m01_axi_awlock),
    .m01_axi_awcache (_if.m01_axi_awcache),
    .m01_axi_awprot (_if.m01_axi_awprot),
    .m01_axi_awqos (_if.m01_axi_awqos),
    .m01_axi_awregion (_if.m01_axi_awregion),
    .m01_axi_awuser (_if.m01_axi_awuser),
    .m01_axi_awvalid (_if.m01_axi_awvalid),
    .m01_axi_awready (_if.m01_axi_awready),
    .m01_axi_wdata (_if.m01_axi_wdata),
    .m01_axi_wstrb (_if.m01_axi_wstrb),
    .m01_axi_wlast (_if.m01_axi_wlast),
    .m01_axi_wuser (_if.m01_axi_wuser),
    .m01_axi_wvalid (_if.m01_axi_wvalid),
    .m01_axi_wready (_if.m01_axi_wready),
    .m01_axi_bid (_if.m01_axi_bid),
    .m01_axi_bresp (_if.m01_axi_bresp),
    .m01_axi_buser (_if.m01_axi_buser),
    .m01_axi_bvalid (_if.m01_axi_bvalid),
    .m01_axi_bready (_if.m01_axi_bready),
    .m01_axi_arid (_if.m01_axi_arid),
    .m01_axi_araddr (_if.m01_axi_araddr),
    .m01_axi_arlen (_if.m01_axi_arlen),
    .m01_axi_arsize (_if.m01_axi_arsize),
    .m01_axi_arburst (_if.m01_axi_arburst),
    .m01_axi_arlock (_if.m01_axi_arlock),
    .m01_axi_arcache (_if.m01_axi_arcache),
    .m01_axi_arprot (_if.m01_axi_arprot),
    .m01_axi_arqos (_if.m01_axi_arqos),
    .m01_axi_arregion (_if.m01_axi_arregion),
    .m01_axi_aruser (_if.m01_axi_aruser),
    .m01_axi_arvalid (_if.m01_axi_arvalid),
    .m01_axi_arready (_if.m01_axi_arready),
    .m01_axi_rid (_if.m01_axi_rid),
    .m01_axi_rdata (_if.m01_axi_rdata),
    .m01_axi_rresp (_if.m01_axi_rresp),
    .m01_axi_rlast (_if.m01_axi_rlast),
    .m01_axi_ruser (_if.m01_axi_ruser),
    .m01_axi_rvalid (_if.m01_axi_rvalid),
    .m01_axi_rready (_if.m01_axi_rready),
  );

endmodule
