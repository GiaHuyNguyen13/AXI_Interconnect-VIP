interface vir_interface (input bit clk);

endinterface