class item extends uvm_sequence_item;
    `uvm_object_utils(item)

endclass                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                