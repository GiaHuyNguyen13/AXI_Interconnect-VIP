interface interface (input bit clk);
    logic rst;

    /*
     * AXI slave interface
     */
    logic [7:0]  s00_axi_awid;        // 8 bits (ID_WIDTH)
    logic [31:0] s00_axi_awaddr;      // 32 bits (ADDR_WIDTH)
    logic [7:0]  s00_axi_awlen;       // 8 bits (fixed)
    logic [2:0]  s00_axi_awsize;      // 3 bits (fixed)
    logic [1:0]  s00_axi_awburst;     // 2 bits (fixed)
    logic        s00_axi_awlock;      // 1 bit (fixed)
    logic [3:0]  s00_axi_awcache;     // 4 bits (fixed)
    logic [2:0]  s00_axi_awprot;      // 3 bits (fixed)
    logic [3:0]  s00_axi_awqos;       // 4 bits (fixed)
    logic [0:0]  s00_axi_awuser;      // 1 bit (AWUSER_WIDTH)
    logic        s00_axi_awvalid;     // 1 bit (fixed)
    logic        s00_axi_awready;     // 1 bit (fixed)
    logic [31:0] s00_axi_wdata;       // 32 bits (DATA_WIDTH)
    logic [3:0]  s00_axi_wstrb;       // 4 bits (STRB_WIDTH)
    logic        s00_axi_wlast;       // 1 bit (fixed)
    logic [0:0]  s00_axi_wuser;       // 1 bit (WUSER_WIDTH)
    logic        s00_axi_wvalid;      // 1 bit (fixed)
    logic        s00_axi_wready;      // 1 bit (fixed)
    logic [7:0]  s00_axi_bid;         // 8 bits (ID_WIDTH)
    logic [1:0]  s00_axi_bresp;       // 2 bits (fixed)
    logic [0:0]  s00_axi_buser;       // 1 bit (BUSER_WIDTH)
    logic        s00_axi_bvalid;      // 1 bit (fixed)
    logic        s00_axi_bready;      // 1 bit (fixed)
    logic [7:0]  s00_axi_arid;        // 8 bits (ID_WIDTH)
    logic [31:0] s00_axi_araddr;      // 32 bits (ADDR_WIDTH)
    logic [7:0]  s00_axi_arlen;       // 8 bits (fixed)
    logic [2:0]  s00_axi_arsize;      // 3 bits (fixed)
    logic [1:0]  s00_axi_arburst;     // 2 bits (fixed)
    logic        s00_axi_arlock;      // 1 bit (fixed)
    logic [3:0]  s00_axi_arcache;     // 4 bits (fixed)
    logic [2:0]  s00_axi_arprot;      // 3 bits (fixed)
    logic [3:0]  s00_axi_arqos;       // 4 bits (fixed)
    logic [0:0]  s00_axi_aruser;      // 1 bit (ARUSER_WIDTH)
    logic        s00_axi_arvalid;     // 1 bit (fixed)
    logic        s00_axi_arready;     // 1 bit (fixed)
    logic [7:0]  s00_axi_rid;         // 8 bits (ID_WIDTH)
    logic [31:0] s00_axi_rdata;       // 32 bits (DATA_WIDTH)
    logic [1:0]  s00_axi_rresp;       // 2 bits (fixed)
    logic        s00_axi_rlast;       // 1 bit (fixed)
    logic [0:0]  s00_axi_ruser;       // 1 bit (RUSER_WIDTH)
    logic        s00_axi_rvalid;      // 1 bit (fixed)
    logic        s00_axi_rready;      // 1 bit (fixed)

    logic [7:0]  s01_axi_awid;        // 8 bits (ID_WIDTH)
    logic [31:0] s01_axi_awaddr;      // 32 bits (ADDR_WIDTH)
    logic [7:0]  s01_axi_awlen;       // 8 bits (fixed)
    logic [2:0]  s01_axi_awsize;      // 3 bits (fixed)
    logic [1:0]  s01_axi_awburst;     // 2 bits (fixed)
    logic        s01_axi_awlock;      // 1 bit (fixed)
    logic [3:0]  s01_axi_awcache;     // 4 bits (fixed)
    logic [2:0]  s01_axi_awprot;      // 3 bits (fixed)
    logic [3:0]  s01_axi_awqos;       // 4 bits (fixed)
    logic [0:0]  s01_axi_awuser;      // 1 bit (AWUSER_WIDTH)
    logic        s01_axi_awvalid;     // 1 bit (fixed)
    logic        s01_axi_awready;     // 1 bit (fixed)
    logic [31:0] s01_axi_wdata;       // 32 bits (DATA_WIDTH)
    logic [3:0]  s01_axi_wstrb;       // 4 bits (STRB_WIDTH)
    logic        s01_axi_wlast;       // 1 bit (fixed)
    logic [0:0]  s01_axi_wuser;       // 1 bit (WUSER_WIDTH)
    logic        s01_axi_wvalid;      // 1 bit (fixed)
    logic        s01_axi_wready;      // 1 bit (fixed)
    logic [7:0]  s01_axi_bid;         // 8 bits (ID_WIDTH)
    logic [1:0]  s01_axi_bresp;       // 2 bits (fixed)
    logic [0:0]  s01_axi_buser;       // 1 bit (BUSER_WIDTH)
    logic        s01_axi_bvalid;      // 1 bit (fixed)
    logic        s01_axi_bready;      // 1 bit (fixed)
    logic [7:0]  s01_axi_arid;        // 8 bits (ID_WIDTH)
    logic [31:0] s01_axi_araddr;      // 32 bits (ADDR_WIDTH)
    logic [7:0]  s01_axi_arlen;       // 8 bits (fixed)
    logic [2:0]  s01_axi_arsize;      // 3 bits (fixed)
    logic [1:0]  s01_axi_arburst;     // 2 bits (fixed)
    logic        s01_axi_arlock;      // 1 bit (fixed)
    logic [3:0]  s01_axi_arcache;     // 4 bits (fixed)
    logic [2:0]  s01_axi_arprot;      // 3 bits (fixed)
    logic [3:0]  s01_axi_arqos;       // 4 bits (fixed)
    logic [0:0]  s01_axi_aruser;      // 1 bit (ARUSER_WIDTH)
    logic        s01_axi_arvalid;     // 1 bit (fixed)
    logic        s01_axi_arready;     // 1 bit (fixed)
    logic [7:0]  s01_axi_rid;         // 8 bits (ID_WIDTH)
    logic [31:0] s01_axi_rdata;       // 32 bits (DATA_WIDTH)
    logic [1:0]  s01_axi_rresp;       // 2 bits (fixed)
    logic        s01_axi_rlast;       // 1 bit (fixed)
    logic [0:0]  s01_axi_ruser;       // 1 bit (RUSER_WIDTH)
    logic        s01_axi_rvalid;      // 1 bit (fixed)
    logic        s01_axi_rready;      // 1 bit (fixed)

    /*
     * AXI master interface
     */
    logic [7:0]  m00_axi_awid;        // 8 bits (ID_WIDTH)
    logic [31:0] m00_axi_awaddr;      // 32 bits (ADDR_WIDTH)
    logic [7:0]  m00_axi_awlen;       // 8 bits (fixed)
    logic [2:0]  m00_axi_awsize;      // 3 bits (fixed)
    logic [1:0]  m00_axi_awburst;     // 2 bits (fixed)
    logic        m00_axi_awlock;      // 1 bit (fixed)
    logic [3:0]  m00_axi_awcache;     // 4 bits (fixed)
    logic [2:0]  m00_axi_awprot;      // 3 bits (fixed)
    logic [3:0]  m00_axi_awqos;       // 4 bits (fixed)
    logic [3:0]  m00_axi_awregion;    // 4 bits (fixed)
    logic [0:0]  m00_axi_awuser;      // 1 bit (AWUSER_WIDTH)
    logic        m00_axi_awvalid;     // 1 bit (fixed)
    logic        m00_axi_awready;     // 1 bit (fixed)
    logic [31:0] m00_axi_wdata;       // 32 bits (DATA_WIDTH)
    logic [3:0]  m00_axi_wstrb;       // 4 bits (STRB_WIDTH)
    logic        m00_axi_wlast;       // 1 bit (fixed)
    logic [0:0]  m00_axi_wuser;       // 1 bit (WUSER_WIDTH)
    logic        m00_axi_wvalid;      // 1 bit (fixed)
    logic        m00_axi_wready;      // 1 bit (fixed)
    logic [7:0]  m00_axi_bid;         // 8 bits (ID_WIDTH)
    logic [1:0]  m00_axi_bresp;       // 2 bits (fixed)
    logic [0:0]  m00_axi_buser;       // 1 bit (BUSER_WIDTH)
    logic        m00_axi_bvalid;      // 1 bit (fixed)
    logic        m00_axi_bready;      // 1 bit (fixed)
    logic [7:0]  m00_axi_arid;        // 8 bits (ID_WIDTH)
    logic [31:0] m00_axi_araddr;      // 32 bits (ADDR_WIDTH)
    logic [7:0]  m00_axi_arlen;       // 8 bits (fixed)
    logic [2:0]  m00_axi_arsize;      // 3 bits (fixed)
    logic [1:0]  m00_axi_arburst;     // 2 bits (fixed)
    logic        m00_axi_arlock;      // 1 bit (fixed)
    logic [3:0]  m00_axi_arcache;     // 4 bits (fixed)
    logic [2:0]  m00_axi_arprot;      // 3 bits (fixed)
    logic [3:0]  m00_axi_arqos;       // 4 bits (fixed)
    logic [3:0]  m00_axi_arregion;    // 4 bits (fixed)
    logic [0:0]  m00_axi_aruser;      // 1 bit (ARUSER_WIDTH)
    logic        m00_axi_arvalid;     // 1 bit (fixed)
    logic        m00_axi_arready;     // 1 bit (fixed)
    logic [7:0]  m00_axi_rid;         // 8 bits (ID_WIDTH)
    logic [31:0] m00_axi_rdata;       // 32 bits (DATA_WIDTH)
    logic [1:0]  m00_axi_rresp;       // 2 bits (fixed)
    logic        m00_axi_rlast;       // 1 bit (fixed)
    logic [0:0]  m00_axi_ruser;       // 1 bit (RUSER_WIDTH)
    logic        m00_axi_rvalid;      // 1 bit (fixed)
    logic        m00_axi_rready;      // 1 bit (fixed)


    logic [7:0]  m01_axi_awid;        // 8 bits (ID_WIDTH)
    logic [31:0] m01_axi_awaddr;      // 32 bits (ADDR_WIDTH)
    logic [7:0]  m01_axi_awlen;       // 8 bits (fixed)
    logic [2:0]  m01_axi_awsize;      // 3 bits (fixed)
    logic [1:0]  m01_axi_awburst;     // 2 bits (fixed)
    logic        m01_axi_awlock;      // 1 bit (fixed)
    logic [3:0]  m01_axi_awcache;     // 4 bits (fixed)
    logic [2:0]  m01_axi_awprot;      // 3 bits (fixed)
    logic [3:0]  m01_axi_awqos;       // 4 bits (fixed)
    logic [3:0]  m01_axi_awregion;    // 4 bits (fixed)
    logic [0:0]  m01_axi_awuser;      // 1 bit (AWUSER_WIDTH)
    logic        m01_axi_awvalid;     // 1 bit (fixed)
    logic        m01_axi_awready;     // 1 bit (fixed)
    logic [31:0] m01_axi_wdata;       // 32 bits (DATA_WIDTH)
    logic [3:0]  m01_axi_wstrb;       // 4 bits (STRB_WIDTH)
    logic        m01_axi_wlast;       // 1 bit (fixed)
    logic [0:0]  m01_axi_wuser;       // 1 bit (WUSER_WIDTH)
    logic        m01_axi_wvalid;      // 1 bit (fixed)
    logic        m01_axi_wready;      // 1 bit (fixed)
    logic [7:0]  m01_axi_bid;         // 8 bits (ID_WIDTH)
    logic [1:0]  m01_axi_bresp;       // 2 bits (fixed)
    logic [0:0]  m01_axi_buser;       // 1 bit (BUSER_WIDTH)
    logic        m01_axi_bvalid;      // 1 bit (fixed)
    logic        m01_axi_bready;      // 1 bit (fixed)
    logic [7:0]  m01_axi_arid;        // 8 bits (ID_WIDTH)
    logic [31:0] m01_axi_araddr;      // 32 bits (ADDR_WIDTH)
    logic [7:0]  m01_axi_arlen;       // 8 bits (fixed)
    logic [2:0]  m01_axi_arsize;      // 3 bits (fixed)
    logic [1:0]  m01_axi_arburst;     // 2 bits (fixed)
    logic        m01_axi_arlock;      // 1 bit (fixed)
    logic [3:0]  m01_axi_arcache;     // 4 bits (fixed)
    logic [2:0]  m01_axi_arprot;      // 3 bits (fixed)
    logic [3:0]  m01_axi_arqos;       // 4 bits (fixed)
    logic [3:0]  m01_axi_arregion;    // 4 bits (fixed)
    logic [0:0]  m01_axi_aruser;      // 1 bit (ARUSER_WIDTH)
    logic        m01_axi_arvalid;     // 1 bit (fixed)
    logic        m01_axi_arready;     // 1 bit (fixed)
    logic [7:0]  m01_axi_rid;         // 8 bits (ID_WIDTH)
    logic [31:0] m01_axi_rdata;       // 32 bits (DATA_WIDTH)
    logic [1:0]  m01_axi_rresp;       // 2 bits (fixed)
    logic        m01_axi_rlast;       // 1 bit (fixed)
    logic [0:0]  m01_axi_ruser;       // 1 bit (RUSER_WIDTH)
    logic        m01_axi_rvalid;      // 1 bit (fixed)
    logic        m01_axi_rready;      // 1 bit (fixed)

endinterface